/*******************
*     a1a1 a2a2
*    f h  i  j b
*    f  h i j  b
*     g1g1 g2g2
*    e  m l k  c
*    e m  l  k c
*     d1d1 d2d2
*
*  FEDCBA9876543210
*  aabcddefgghijklm
*  12  12  12
*******************/
module charROM(
input wire [7:0] ascii,
output wire [15:0] segments
);

reg [15:0] seg;

assign segments[15:0] = seg [15:0];

always 
begin
	case(ascii)
		"0": seg = 16'b0000000011111111;
		"1": seg = 16'b1100111111110111;
		"2": seg = 16'b0001000100111111;
		"3": seg = 16'b0000001110111111;
		"4": seg = 16'b1100111000111111;
		"5": seg = 16'b0010001000111111;
		"6": seg = 16'b0010000000111111;
		"7": seg = 16'b0000111111111111;
		"8": seg = 16'b0000000000111111;
		"9": seg = 16'b0000111000111111;
		":": seg = 16'b1111111111101101;
		";": seg = 16'b1111111111101110;
		"<": seg = 16'b1111111111110011;
		"=": seg = 16'b1111001100111111;
		">": seg = 16'b1111111111011110;
		"?": seg = 16'b0001111110111101;
		"@": seg = 16'b0001000010110111;
		"A": seg = 16'b0000110000111111;
		"B": seg = 16'b0000001110101101;
		"C": seg = 16'b0011000011111111;
		"D": seg = 16'b0000001111101101;
		"E": seg = 16'b0011000000111111;
		"F": seg = 16'b0011110001111111;
		"G": seg = 16'b0010000010111111;
		"H": seg = 16'b1100110000111111;
		"I": seg = 16'b1111111111101101;
		"J": seg = 16'b1100000111111111;
		"K": seg = 16'b1111110011110011;
		"L": seg = 16'b1111000011111111;
		"M": seg = 16'b1100110011010111;
		"N": seg = 16'b1100110011011011;
		"O": seg = 16'b0000000011111111;
		"P": seg = 16'b0001110000111111;
		"Q": seg = 16'b0000000011111011;
		"R": seg = 16'b0001110000111011;
		"S": seg = 16'b0010001110011111;
		"T": seg = 16'b0011111111101101;
		"U": seg = 16'b1100000011111111;
		"V": seg = 16'b1111110011110110;
		"W": seg = 16'b1100110011111010;
		"X": seg = 16'b1111111111010010;
		"Y": seg = 16'b1111111111010101;
		"Z": seg = 16'b0011001111110110;
		"[": seg = 16'b0111010011111111;
		"\\": seg = 16'b1111111111011110;
		"]": seg = 16'b1000101111111111;
		"^": seg = 16'b1111111011011111;
		"_": seg = 16'b1111001111111111;
		"`": seg = 16'b1111111111011111;

		default : seg = 16'b1111111111111111;
	endcase
end //always

endmodule
